

package INSTRUCTION_FETCH_PKG;

endpackage